module PS2(
	input wire clk,
	input wire reset_n,
	
	// RISC-V interface
	input  wire [ 9:0] r_addr,
	input  wire [31:0] r_din,
	output reg  [31:0] r_dout,
	input  wire [ 3:0] r_lane,
	input  wire        r_wr,
	input  wire        r_valid,
	output reg         r_ready,

	// CPU interface
	input wire [11:0] port,
	output reg [7:0] dout,
	input wire [7:0] din,
	input wire cpu_iordin,
	output reg cpu_iordout,
	input wire cpu_iowrin,
	output reg cpu_iowrout,

	output reg irq1
);

reg   [7:0] buffer [0:15];
reg   [3:0] rp;
reg   [3:0] wp;
reg   [4:0] count;

wire iord = cpu_iordout ^ cpu_iordin;
wire iowr = cpu_iowrout ^ cpu_iowrin;

reg cs_60h;
reg cs_61h;

always @(negedge clk)
begin
	cs_60h <= port == 12'h060;
	cs_61h <= port == 12'h061;
end

wire [3:0] wp_next;
assign wp_next = wp + 1'd1;

always @(posedge clk)
begin
	cpu_iordout <= cpu_iordin;
	cpu_iowrout <= cpu_iowrin;
	
	dout <= buffer[rp];
	irq1 <= rp != wp;

	r_ready <= 1'b0;
	
	if (cs_61h && iowr)
	begin
		if (rp != wp)
			rp <= rp + 1'd1;
	end
	else if (r_valid)
	begin
		r_ready <= 1'b1;
		if (r_valid & ~r_ready)
		begin
			if (wp_next != rp)
			begin
				buffer[wp] <= r_din[7:0];
				wp <= wp + 1'd1;
			end
		end
	end
end

endmodule
